/*
 * Ultra wide range test
*/

`define WIDTH 256
`define operator not
`include "../generic/replicate_any_width_unary_test.v"