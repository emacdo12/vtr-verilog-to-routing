/*
 * Wide range test
*/

`define WIDTH 3
`define operator not
`include "../generic/replicate_any_width_unary_test.v"