/*
 * Integer wide range test
*/

`define WIDTH 32
`define operator and
`include "../generic/range_any_width_binary_test.v"