/*
 * Wide range test
*/

`define WIDTH 3
`define operator or
`include "../generic/range_any_width_binary_test.v"