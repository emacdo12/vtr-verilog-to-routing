`define WIDTH 3 

module simple_op(input in,output out);
	assign out = in;
endmodule 