/*
 * Integer wide range test
*/

`define WIDTH 32
`define operator not
`include "../generic/range_any_width_unary_test.v"