/*
 * Wide range test
*/

`define WIDTH 3
`define operator xor
`include "../generic/range_any_width_binary_test.v"