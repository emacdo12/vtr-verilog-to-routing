`define BINARY_OP(out,a,b) or(out, a, b);
`include "../generic/wire_test.v"