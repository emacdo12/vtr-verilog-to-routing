/*
 * Wide range test
*/

`define WIDTH 3
`define operator buf
`include "../generic/range_any_width_unary_test.v"