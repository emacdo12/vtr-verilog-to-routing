/*
 * Wide range test
*/

`define WIDTH 3
`define operator buf
`include "../generic/replicate_any_width_unary_test.v"