`define UNARY_OP(out,a) not(out, a);
`include "../generic/wire_test.v"