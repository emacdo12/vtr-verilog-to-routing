`define BINARY_OP(out,a,b) nor(out, a, b);
`include "../generic/wire_test.v"