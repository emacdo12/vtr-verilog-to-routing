module simple_op(a,b,c);
input a;
input b;

output c;

wire a,b,c;

assign c = a&b;

endmodule