/*
 * Integer wide range test
*/

`define WIDTH 32
`define operator buf
`include "../generic/range_any_width_unary_test.v"