`define BINARY_OP(out,a,b) xor(out, a, b);
`include "../generic/wire_test.v"