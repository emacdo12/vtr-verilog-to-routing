`define BINARY_OP(out,a,b) and(out, a, b);
`include "../generic/wire_test.v"