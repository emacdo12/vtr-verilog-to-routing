/*
 * Integer wide range test
*/

`define WIDTH 32
`define operator xor
`include "../generic/replicate_any_width_binary_test.v"