/*
 * Integer wide range test
*/

`define WIDTH 32
`define operator xnor
`include "../generic/range_any_width_binary_test.v"